i am in fourth 
fourth file change
