i am in vineet branch
in vineet 
