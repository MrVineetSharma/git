i am in third file
